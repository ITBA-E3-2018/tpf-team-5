`include "ImageDrawer.v"
//Modulo que se encarga de verficar que ImageDrawer dibuja
//exitosamente los simbolos en la pantalla.
module ImageDrawer_tb;

 ImageDrawer inst(hours,minutes,seconds,milliseconds,enable,row,column,r,g,b);


endmodule // ImageDrawer_tb